module winograd(inp10, inp11, inp12, inp13 ,inp20,inp21,inp22,inp23,inp30,inp31,
inp32,inp33,inp40,inp41,inp42,inp43,ker10,ker11,ker12,ker20,ker21,ker22,
ker30,ker31,ker32,out10,out11,out20,out21);

input [7:0] inp10, inp11, inp12, inp13;
input [7:0] inp20, inp21, inp22, inp23;
input [7:0] inp30, inp31, inp32, inp33;
input [7:0] inp40, inp41, inp42, inp43;

input [7:0] ker10, ker11, ker12;
input [7:0] ker20, ker21, ker22;
input [7:0] ker30, ker31, ker32;

output reg [7:0] out10,out11;
output reg [7:0] out20,out21;

reg [7:0] pre1 [1:0];
reg [7:0] pre2 [1:0];

reg [7:0] pre_out1 [1:0];
reg [7:0] pre_out2 [1:0];

reg [7:0] p1 [2:0];
reg [7:0] p2 [2:0];
reg [7:0] p3 [2:0];
reg [7:0] p4 [2:0];

reg [7:0] q1 [3:0];
reg [7:0] q2 [3:0];
reg [7:0] q3 [3:0];
reg [7:0] q4 [3:0];

reg [7:0] s1 [3:0];
reg [7:0] s2 [3:0];
reg [7:0] s3 [3:0];
reg [7:0] s4 [3:0];

reg [7:0] t1 [3:0];
reg [7:0] t2 [3:0];
reg [7:0] t3 [3:0];
reg [7:0] t4 [3:0];

reg [7:0] qt1 [3:0];
reg [7:0] qt2 [3:0];
reg [7:0] qt3 [3:0];
reg [7:0] qt4 [3:0];

reg [7:0] y1 [3:0];
reg [7:0] y2 [3:0];

//reg [7:0] a1 [1:0] = {8'h01, 8'h00}; // a1 = [1, 0]
//reg [7:0] a2 [1:0] = {8'h01, 8'h01}; // a2 = [1, 1]
//reg [7:0] a3 [1:0] = {8'h01, 8'hFF}; // a3 = [1, -1]
//reg [7:0] a4 [1:0] = {8'h00, 8'hFF}; // a4 = [0, -1]

//reg [7:0] b1 [3:0]  = {8'h01, 8'h00, 8'hFF, 8'h00}; // b1 = [1, 0, -1, 0]
//reg [7:0] b2 [3:0]  = {8'h00, 8'h01, 8'h01, 8'h00}; // b2 = [0, 1, 1, 0]
//reg [7:0] b3 [3:0]  = {8'h00, 8'hFF, 8'h01, 8'h00}; // b3 = [0,-1, 1, 0]
//reg [7:0] b4 [3:0]  = {8'h00, 8'h01, 8'h00, 8'hFF}; // b4 = [0, 1, 0, -1]

//reg [7:0] bT1 [3:0]  = {8'h01, 8'h00, 8'h00, 8'h00}; // b1 = [1, 0, 0, 0]
//reg [7:0] bT2 [3:0]  = {8'h00, 8'h01, 8'hFF, 8'h01}; // b2 = [0, 1, -1, 1]
//reg [7:0] bT3 [3:0]  = {8'hFF, 8'h01, 8'h01, 8'h00}; // b3 = [-1, 1, 1, 0]
//reg [7:0] bT4 [3:0]  = {8'h00, 8'h00, 8'h00, 8'hFF}; // b4 = [0, 0, 0, -1]

//reg [7:0] g1 [2:0] = {8'h02, 8'h00, 8'h00}; // g1 = [2, 0, 0]
//reg [7:0] g2 [2:0] = {8'h01, 8'h01, 8'h01}; // g2 = [1, 1, 1]
//reg [7:0] g3 [2:0] = {8'h01, 8'hFF, 8'h01}; // g3 = [1, -1, 1]
//reg [7:0] g4 [2:0] = {8'h00, 8'h00, 8'h02}; // g4 = [0, 0, 2]

//reg [7:0] gT1 [3:0] = {8'h02, 8'h01, 8'h01, 8'h00}; // g1 = [2, 1, 1 , 0]
//reg [7:0] gT2 [3:0] = {8'h00, 8'h01, 8'hFF, 8'h00}; // g2 = [0, 1, -1, 0]
//reg [7:0] gT3 [3:0] = {8'h00, 8'h01, 8'h01, 8'h02}; // g3 = [0, 1, 1, 2]

//reg [7:0] aT1 [3:0] = {8'h01, 8'h01, 8'h01, 8'h00}; // a1 = [1, 1, 1, 0]
//reg [7:0] aT2 [3:0] = {8'h00, 8'h01, 8'hFF, 8'hFF}; // a2 = [0, 1, -1, -1]


reg [7:0] a1 [1:0];
reg [7:0] a2 [1:0];
reg [7:0] a3 [1:0];
reg [7:0] a4 [1:0];

initial begin
    a1[1] = 8'h01;
    a1[0] = 8'h00;
    
    a2[1] = 8'h01;
    a2[0] = 8'h01;
    
    a3[1] = 8'h01;
    a3[0] = 8'hFF;
    
    a4[1] = 8'h00;
    a4[0] = 8'hFF;
end

reg [7:0] bT1 [3:0];
reg [7:0] bT2 [3:0];
reg [7:0] bT3 [3:0];
reg [7:0] bT4 [3:0];

initial begin
    bT1[3] = 8'h01;
    bT1[2] = 8'h00;
    bT1[1] = 8'hFF;
    bT1[0] = 8'h00;
    
    bT2[3] = 8'h00;
    bT2[2] = 8'h01;
    bT2[1] = 8'h01;
    bT2[0] = 8'h00;
    
    bT3[3] = 8'h00;
    bT3[2] = 8'hFF;
    bT3[1] = 8'h01;
    bT3[0] = 8'h00;
    
    bT4[3] = 8'h00;
    bT4[2] = 8'h01;
    bT4[1] = 8'h00;
    bT4[0] = 8'hFF;
end

reg [7:0] b1 [3:0];
reg [7:0] b2 [3:0];
reg [7:0] b3 [3:0];
reg [7:0] b4 [3:0];

initial begin
    b1[3] = 8'h01;
    b1[2] = 8'h00;
    b1[1] = 8'h00;
    b1[0] = 8'h00;
    
    b2[3] = 8'h00;
    b2[2] = 8'h01;
    b2[1] = 8'hFF;
    b2[0] = 8'h01;
    
    b3[3] = 8'hFF;
    b3[2] = 8'h01;
    b3[1] = 8'h01;
    b3[0] = 8'h00;
    
    b4[3] = 8'h00;
    b4[2] = 8'h00;
    b4[1] = 8'h00;
    b4[0] = 8'hFF;
end

reg [7:0] g1 [2:0];
reg [7:0] g2 [2:0];
reg [7:0] g3 [2:0];
reg [7:0] g4 [2:0];

initial begin
    g1[2] = 8'h02;
    g1[1] = 8'h00;
    g1[0] = 8'h00;
    
    g2[2] = 8'h01;
    g2[1] = 8'h01;
    g2[0] = 8'h01;
    
    g3[2] = 8'h01;
    g3[1] = 8'hFF;
    g3[0] = 8'h01;
    
    g4[2] = 8'h00;
    g4[1] = 8'h00;
    g4[0] = 8'h02;
end

reg [7:0] gT1 [3:0];
reg [7:0] gT2 [3:0];
reg [7:0] gT3 [3:0];

initial begin
    gT1[3] = 8'h02;
    gT1[2] = 8'h01;
    gT1[1] = 8'h01;
    gT1[0] = 8'h00;
    
    gT2[3] = 8'h00;
    gT2[2] = 8'h01;
    gT2[1] = 8'hFF;
    gT2[0] = 8'h00;
    
    gT3[3] = 8'h00;
    gT3[2] = 8'h01;
    gT3[1] = 8'h01;
    gT3[0] = 8'h02;
end

reg [7:0] aT1 [3:0];
reg [7:0] aT2 [3:0];

initial begin
    aT1[3] = 8'h01;
    aT1[2] = 8'h01;
    aT1[1] = 8'h01;
    aT1[0] = 8'h00;
    
    aT2[3] = 8'h00;
    aT2[2] = 8'h01;
    aT2[1] = 8'hFF;
    aT2[0] = 8'hFF;
end

reg [7:0] g_gT_multiple = 8'd25; //Its actually decimal 0.25 when 0.5 is taken as common from both G and G transform and multiplied, but its stored as 25 and during operation we can divide it by 100


always @(*)
begin
//G*kernel

//p1[0] = g1[2]*ker10 + g1[1]*ker20 + g1[0]*ker30;
//p1[1] = g1[2]*ker11 + g1[1]*ker21 + g1[0]*ker31;
//p1[2] = g1[2]*ker12 + g1[1]*ker22 + g1[0]*ker32;

//p2[0] = g2[2]*ker10 + g2[1]*ker20 + g2[0]*ker30;
//p2[1] = g2[2]*ker11 + g2[1]*ker21 + g2[0]*ker31;
//p2[2] = g2[2]*ker12 + g2[1]*ker22 + g2[0]*ker32;

//p3[0] = g3[2]*ker10 + g3[1]*ker20 + g3[0]*ker30;
//p3[1] = g3[2]*ker11 + g3[1]*ker21 + g3[0]*ker31;
//p3[2] = g3[2]*ker12 + g3[1]*ker22 + g3[0]*ker32;

//p4[0] = g4[2]*ker10 + g4[1]*ker20 + g4[0]*ker30;
//p4[1] = g4[2]*ker11 + g4[1]*ker21 + g4[0]*ker31;
//p4[2] = g4[2]*ker12 + g4[1]*ker22 + g4[0]*ker32;

p1[2] = g1[2]*ker10 + g1[1]*ker20 + g1[0]*ker30;
p1[1] = g1[2]*ker11 + g1[1]*ker21 + g1[0]*ker31;
p1[0] = g1[2]*ker12 + g1[1]*ker22 + g1[0]*ker32;

p2[2] = g2[2]*ker10 + g2[1]*ker20 + g2[0]*ker30;
p2[1] = g2[2]*ker11 + g2[1]*ker21 + g2[0]*ker31;
p2[0] = g2[2]*ker12 + g2[1]*ker22 + g2[0]*ker32;

p3[2] = g3[2]*ker10 + g3[1]*ker20 + g3[0]*ker30;
p3[1] = g3[2]*ker11 + g3[1]*ker21 + g3[0]*ker31;
p3[0] = g3[2]*ker12 + g3[1]*ker22 + g3[0]*ker32;

p4[2] = g4[2]*ker10 + g4[1]*ker20 + g4[0]*ker30;
p4[1] = g4[2]*ker11 + g4[1]*ker21 + g4[0]*ker31;
p4[0] = g4[2]*ker12 + g4[1]*ker22 + g4[0]*ker32;
   

end


always @(*)
begin
//transformed kernel (G*kernel*GT)
q1[3] = p1[2]*gT1[3] + p1[1]*gT2[3] + p1[0]*gT3[3];
q1[2] = p1[2]*gT1[2] + p1[1]*gT2[2] + p1[0]*gT3[2];
q1[1] = p1[2]*gT1[1] + p1[1]*gT2[1] + p1[0]*gT3[1];
q1[0] = p1[2]*gT1[0] + p1[1]*gT2[0] + p1[0]*gT3[0];

q2[3] = p2[2]*gT1[3] + p2[1]*gT2[3] + p2[0]*gT3[3];
q2[2] = p2[2]*gT1[2] + p2[1]*gT2[2] + p2[0]*gT3[2];
q2[1] = p2[2]*gT1[1] + p2[1]*gT2[1] + p2[0]*gT3[1];
q2[0] = p2[2]*gT1[0] + p2[1]*gT2[0] + p2[0]*gT3[0];

q3[3] = p3[2]*gT1[3] + p3[1]*gT2[3] + p3[0]*gT3[3];
q3[2] = p3[2]*gT1[2] + p3[1]*gT2[2] + p3[0]*gT3[2];
q3[1] = p3[2]*gT1[1] + p3[1]*gT2[1] + p3[0]*gT3[1];
q3[0] = p3[2]*gT1[0] + p3[1]*gT2[0] + p3[0]*gT3[0];

q4[3] = p4[2]*gT1[3] + p4[1]*gT2[3] + p4[0]*gT3[3];
q4[2] = p4[2]*gT1[2] + p4[1]*gT2[2] + p4[0]*gT3[2];
q4[1] = p4[2]*gT1[1] + p4[1]*gT2[1] + p4[0]*gT3[1];
q4[0] = p4[2]*gT1[0] + p4[1]*gT2[0] + p4[0]*gT3[0];


end

always @(*)
begin
//BT*input
s1[3] = bT1[3]*inp10 + bT1[2]*inp20 + bT1[1]*inp30 + bT1[0]*inp40;
s1[2] = bT1[3]*inp11 + bT1[2]*inp21 + bT1[1]*inp31 + bT1[0]*inp41;
s1[1] = bT1[3]*inp12 + bT1[2]*inp22 + bT1[1]*inp32 + bT1[0]*inp42;
s1[0] = bT1[3]*inp13 + bT1[2]*inp23 + bT1[1]*inp33 + bT1[0]*inp43;

s2[3] = bT2[3]*inp10 + bT2[2]*inp20 + bT2[1]*inp30 + bT2[0]*inp40;
s2[2] = bT2[3]*inp11 + bT2[2]*inp21 + bT2[1]*inp31 + bT2[0]*inp41;
s2[1] = bT2[3]*inp12 + bT2[2]*inp22 + bT2[1]*inp32 + bT2[0]*inp42;
s2[0] = bT2[3]*inp13 + bT2[2]*inp23 + bT2[1]*inp33 + bT2[0]*inp43;

s3[3] = bT3[3]*inp10 + bT3[2]*inp20 + bT3[1]*inp30 + bT3[0]*inp40;
s3[2] = bT3[3]*inp11 + bT3[2]*inp21 + bT3[1]*inp31 + bT3[0]*inp41;
s3[1] = bT3[3]*inp12 + bT3[2]*inp22 + bT3[1]*inp32 + bT3[0]*inp42;
s3[0] = bT3[3]*inp13 + bT3[2]*inp23 + bT3[1]*inp33 + bT3[0]*inp43;

s4[3] = bT4[3]*inp10 + bT4[2]*inp20 + bT4[1]*inp30 + bT4[0]*inp40;
s4[2] = bT4[3]*inp11 + bT4[2]*inp21 + bT4[1]*inp31 + bT4[0]*inp41;
s4[1] = bT4[3]*inp12 + bT4[2]*inp22 + bT4[1]*inp32 + bT4[0]*inp42;
s4[0] = bT4[3]*inp13 + bT4[2]*inp23 + bT4[1]*inp33 + bT4[0]*inp43;
end

always @(*)
begin
//transformed feature map (BT*input*B)
t1[3] = s1[3]*b1[3] + s1[2]*b2[3] + s1[1]*b3[3] + s1[0]*b4[3];
t1[2] = s1[3]*b1[2] + s1[2]*b2[2] + s1[1]*b3[2] + s1[0]*b4[2];
t1[1] = s1[3]*b1[1] + s1[2]*b2[1] + s1[1]*b3[1] + s1[0]*b4[1];
t1[0] = s1[3]*b1[0] + s1[2]*b2[0] + s1[1]*b3[0] + s1[0]*b4[0];

t2[3] = s2[3]*b1[3] + s2[2]*b2[3] + s2[1]*b3[3] + s2[0]*b4[3];
t2[2] = s2[3]*b1[2] + s2[2]*b2[2] + s2[1]*b3[2] + s2[0]*b4[2];
t2[1] = s2[3]*b1[1] + s2[2]*b2[1] + s2[1]*b3[1] + s2[0]*b4[1];
t2[0] = s2[3]*b1[0] + s2[2]*b2[0] + s2[1]*b3[0] + s2[0]*b4[0];

t3[3] = s3[3]*b1[3] + s3[2]*b2[3] + s3[1]*b3[3] + s3[0]*b4[3];
t3[2] = s3[3]*b1[2] + s3[2]*b2[2] + s3[1]*b3[2] + s3[0]*b4[2];
t3[1] = s3[3]*b1[1] + s3[2]*b2[1] + s3[1]*b3[1] + s3[0]*b4[1];
t3[0] = s3[3]*b1[0] + s3[2]*b2[0] + s3[1]*b3[0] + s3[0]*b4[0];

t4[3] = s4[3]*b1[3] + s4[2]*b2[3] + s4[1]*b3[3] + s4[0]*b4[3];
t4[2] = s4[3]*b1[2] + s4[2]*b2[2] + s4[1]*b3[2] + s4[0]*b4[2];
t4[1] = s4[3]*b1[1] + s4[2]*b2[1] + s4[1]*b3[1] + s4[0]*b4[1];
t4[0] = s4[3]*b1[0] + s4[2]*b2[0] + s4[1]*b3[0] + s4[0]*b4[0];

end

always @(*)
begin
//Elementwise mult qt
qt1[0] = q1[0]*t1[0];
qt1[1] = q1[1]*t1[1];
qt1[2] = q1[2]*t1[2];
qt1[3] = q1[3]*t1[3];

qt2[0] = q2[0]*t2[0];
qt2[1] = q2[1]*t2[1];
qt2[2] = q2[2]*t2[2];
qt2[3] = q2[3]*t2[3];

qt3[0] = q3[0]*t3[0];
qt3[1] = q3[1]*t3[1];
qt3[2] = q3[2]*t3[2];
qt3[3] = q3[3]*t3[3];

qt4[0] = q4[0]*t4[0];
qt4[1] = q4[1]*t4[1];
qt4[2] = q4[2]*t4[2];
qt4[3] = q4[3]*t4[3];

//AT*QT
y1[3] = aT1[3]*qt1[3] + aT1[2]*qt2[3] + aT1[1]*qt3[3] + aT1[0]*qt4[3];
y1[2] = aT1[3]*qt1[2] + aT1[2]*qt2[2] + aT1[1]*qt3[2] + aT1[0]*qt4[2];
y1[1] = aT1[3]*qt1[1] + aT1[2]*qt2[1] + aT1[1]*qt3[1] + aT1[0]*qt4[1];
y1[0] = aT1[3]*qt1[0] + aT1[2]*qt2[0] + aT1[1]*qt3[0] + aT1[0]*qt4[0];

y2[3] = aT2[3]*qt1[3] + aT2[2]*qt2[3] + aT2[1]*qt3[3] + aT2[0]*qt4[3];
y2[2] = aT2[3]*qt1[2] + aT2[2]*qt2[2] + aT2[1]*qt3[2] + aT2[0]*qt4[2];
y2[1] = aT2[3]*qt1[1] + aT2[2]*qt2[1] + aT2[1]*qt3[1] + aT2[0]*qt4[1];
y2[0] = aT2[3]*qt1[0] + aT2[2]*qt2[0] + aT2[1]*qt3[0] + aT2[0]*qt4[0];

//AT*QT*A - Output Transformation
pre_out1[1] = y1[3]*a1[1] + y1[2]*a2[1] + y1[1]*a3[1] + y1[0]*a4[1];
pre_out1[0] = y1[3]*a1[0] + y1[2]*a2[0] + y1[1]*a3[0] + y1[0]*a4[0];

pre_out2[1] = y2[3]*a1[1] + y2[2]*a2[1] + y2[1]*a3[1] + y2[0]*a4[1];
pre_out2[0] = y2[3]*a1[0] + y2[2]*a2[0] + y2[1]*a3[0] + y2[0]*a4[0];

pre1[1] = pre_out1[1]/4;
pre1[0] = pre_out1[0]/4;

pre2[1] = pre_out2[1]/4;
pre2[0] = pre_out2[0]/4;
 
 out10 = (pre1[1][5] == 1'b1)? {2'b11,pre1[1][5:0]} : (pre1[1]);
 out11 = (pre1[0][5] == 1'b1)? {2'b11,pre1[0][5:0]} : (pre1[0]);
 
  out20 = (pre2[1][5] == 1'b1)? {2'b11,pre2[1][5:0]} : (pre2[1]);
  out21 = (pre2[0][5] == 1'b1)? {2'b11,pre2[0][5:0]} : (pre2[0]);


end


endmodule