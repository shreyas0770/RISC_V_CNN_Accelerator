module and_gate(a,b,out);
input a,b,c;
output out;

assign out = a & b;
endmodule
