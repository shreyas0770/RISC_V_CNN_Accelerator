module and_gate(a,b,y);
input a,b,c;
output y;

assign y = a & b;
endmodule
